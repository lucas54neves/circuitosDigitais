entity decodificador is
port(
    signed_int: IN BIT_VECTOR(4 DOWNTO 0);
    digits: OUT BIT_VECTOR(13 DOWNTO 0));
end decodificador;
 
architecture behavioral of decodificador is
begin
    WITH signed_int SELECT
                     
        digits <=
            -- Positive values:
            NOT("11111101111110") WHEN "00000", -- 00
            NOT("11111100110000") WHEN "00001", -- 01
            NOT("11111101101101") WHEN "00010", -- 02
            NOT("11111101111001") WHEN "00011", -- 03
            NOT("11111100110011") WHEN "00100", -- 04
            NOT("11111101011011") WHEN "00101", -- 05
            NOT("11111101011111") WHEN "00110", -- 06
            NOT("11111101110000") WHEN "00111", -- 07
            NOT("11111101111111") WHEN "01000", -- 08
            NOT("11111101110011") WHEN "01001", -- 09
            NOT("01100001111110") WHEN "01010", -- 10
            NOT("01100000110000") WHEN "01011", -- 11
            NOT("01100001101101") WHEN "01100", -- 12
            NOT("01100001111001") WHEN "01101", -- 13
            NOT("01100000110011") WHEN "01110", -- 14     
            NOT("01100001011011") WHEN "01111", -- 15
            NOT("01100001011111") WHEN "10000", -- 16
            NOT("01100001110000") WHEN "10001", -- 17
            NOT("01100001111111") WHEN "10010", -- 18
            NOT("01100001110011") WHEN "10011", -- 19
            NOT("11011011111110") WHEN "10100", -- 20
            NOT("11011010110000") WHEN "10101", -- 21
            NOT("11011011101101") WHEN "10110", -- 22
            NOT("11011011111001") WHEN "10111", -- 23
            NOT("11011010110011") WHEN "11000", -- 24
            NOT("11011011011011") WHEN "11001", -- 25
            NOT("11011011011111") WHEN "11010", -- 26
            NOT("11011011110000") WHEN "11011", -- 27
            NOT("11011011111111") WHEN "11100", -- 28
            NOT("11011011110011") WHEN "11101", -- 29
            NOT("11110011111110") WHEN "11110", -- 30    
            NOT("11110010110000") WHEN "11111"; -- 31
                 
end behavioral;